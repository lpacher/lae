//
// Behavioural implementation of a 5-bit/32-bit one-hot decoder using a for-loop statement.
//
// Luca Pacher - pacher@to.infn.it
// Spring 2020
//


`timescale 1ns / 100ps

module OneHotDecoder (

   input  wire [4:0]  Bin,      //  5-bit base-2 binary input code
   output reg  [31:0] Bout      // 32-bit one-hot output code
 
   ) ;

/*
   always @(*) begin

      case (Bin)

         5'b00000 : Bout = 32'b00000000000000000000000000000001 ;
         5'b00001 : Bout = 32'b00000000000000000000000000000010 ;
         5'b00010 : Bout = 32'b00000000000000000000000000000100 ;
         5'b00011 : Bout = 32'b00000000000000000000000000001000 ;
         5'b00100 : Bout = 32'b00000000000000000000000000010000 ;
         5'b00101 : Bout = 32'b00000000000000000000000000100000 ;
         5'b00110 : Bout = 32'b00000000000000000000000001000000 ;
         5'b00111 : Bout = 32'b00000000000000000000000010000000 ;
         5'b01000 : Bout = 32'b00000000000000000000000100000000 ;
         5'b01001 : Bout = 32'b00000000000000000000001000000000 ;
         5'b01010 : Bout = 32'b00000000000000000000010000000000 ;
         5'b01011 : Bout = 32'b00000000000000000000100000000000 ;
         5'b01100 : Bout = 32'b00000000000000000001000000000000 ;
         5'b01101 : Bout = 32'b00000000000000000010000000000000 ;
         5'b01110 : Bout = 32'b00000000000000000100000000000000 ;
         5'b01111 : Bout = 32'b00000000000000001000000000000000 ;
         5'b10000 : Bout = 32'b00000000000000010000000000000000 ;
         5'b10001 : Bout = 32'b00000000000000100000000000000000 ;
         5'b10010 : Bout = 32'b00000000000001000000000000000000 ;
         5'b10011 : Bout = 32'b00000000000010000000000000000000 ;
         5'b10100 : Bout = 32'b00000000000100000000000000000000 ;
         5'b10101 : Bout = 32'b00000000001000000000000000000000 ;
         5'b10110 : Bout = 32'b00000000010000000000000000000000 ;
         5'b10111 : Bout = 32'b00000000100000000000000000000000 ;
         5'b11000 : Bout = 32'b00000001000000000000000000000000 ;
         5'b11001 : Bout = 32'b00000010000000000000000000000000 ;
         5'b11010 : Bout = 32'b00000100000000000000000000000000 ;
         5'b11011 : Bout = 32'b00001000000000000000000000000000 ;
         5'b11100 : Bout = 32'b00010000000000000000000000000000 ;
         5'b11101 : Bout = 32'b00100000000000000000000000000000 ;
         5'b11110 : Bout = 32'b01000000000000000000000000000000 ;
         5'b11111 : Bout = 32'b10000000000000000000000000000000 ;

         default  : Bout = 32'b00000000000000000000000000000001 ;

      endcase
   end   // always
*/

   integer i ;

   always @(*) begin

      for(i=0; i < 32; i=i+1) begin

         Bout[i] = (Bin[4:0] ==i) ;      // this is equivalent to (Bin[4:0] == i) ? 1'b1 : 1'b0 ;

         //if (Bin[4:0] == i) begin
         //   Bout[i] = 1'b1 ;
         //end
         //else begin 
         //   Bout[i] = 1'b0 ;
         //end

      end  // for
   end  // always

endmodule

